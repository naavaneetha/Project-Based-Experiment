library verilog;
use verilog.vl_types.all;
entity projectbased_vlg_check_tst is
    port(
        G1              : in     vl_logic;
        G2              : in     vl_logic;
        G3              : in     vl_logic;
        PG              : in     vl_logic;
        PR              : in     vl_logic;
        R1              : in     vl_logic;
        R2              : in     vl_logic;
        R3              : in     vl_logic;
        Y1              : in     vl_logic;
        Y2              : in     vl_logic;
        Y3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end projectbased_vlg_check_tst;
