library verilog;
use verilog.vl_types.all;
entity projectbased_vlg_vec_tst is
end projectbased_vlg_vec_tst;
